library verilog;
use verilog.vl_types.all;
entity down_counter_testbench is
end down_counter_testbench;
