library verilog;
use verilog.vl_types.all;
entity johnson_counter_testbench is
end johnson_counter_testbench;
